module test(input a,b,output out1,out2);
assign out1 = a&b;
assign out2 = a|b;
endmodule